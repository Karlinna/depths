[PLAYER]
Name:Anna
LocX:6
LocY:1
Class:WARRIOR
Gender:FEMALE
Image:C:/Users/IBM_ADMIN/source/repos/depths2/Depths/bin/Debug/depths_images/female/human_female_warrior.gif
Level:1
Exp:0
[PLAYER]
[STORY]
[DIALOGUE]
Test:"You are at 3, 1, warrior."
[DIALOGUE]
[DIALOGUE]
Test:"This is where you engage a battle, Anna."
[DIALOGUE]
[DIALOGUE]
Anna:"You wanted this, Test."
[DIALOGUE]
[DIALOGUE]
Anna:"This is a shallow speak at 9,5"
[DIALOGUE]
[DIALOGUE]
Narrator:"This is narration at 9,5"
[DIALOGUE]
[DIALOGUE]
Anna:"Shallow speak with only player speech."
[DIALOGUE]
[DIALOGUE]
Anna:"Should it cause error if no narrator?"
[DIALOGUE]
[DIALOGUE]
Anna:"Probably not."
[DIALOGUE]
[DIALOGUE]
Narrator:"Lady and Lady"
[DIALOGUE]
[MAPCONDITION]
exists:False
startIndex:0
endIndex:2
[ENEMY]
name:Test
LocX:3
LocY:1
[ENEMY]
[MAPCONDITION]
[MAPCONDITION]
exists:True
startIndex:3
endIndex:4
[NARRATOR]
name:Narrator
LocX:9
LocY:5
[NARRATOR]
[MAPCONDITION]
[MAPCONDITION]
exists:True
startIndex:5
endIndex:8
[NARRATOR]
name:Narrator
LocX:9
LocY:6
[NARRATOR]
[MAPCONDITION]
[STORY]
